module lab5_tb;
reg [31:0] x, y;
wire [31:0] r;

lab5 uut(r, x, y);

initial
begin
	//x[31] = 1'b0; x[30:23] = 8'b0000_0000; x[22:0] = 23'b000_0000_0000_0000_0000_0000;
	//y[31] = 1'b0; y[30:23] = 8'b0000_0000; y[22:0] = 23'b000_0000_0000_0000_0000_0000;
	
	x = 32'b00111111100100000000000000000000; //1.125
	y = 32'b01000000011000000000000000000000; //3.5
	//r = 01000000011111000000000000000000 = 3.9375
	
	//x = 32'b00000000000000000000000000000011;
	//y = 32'b00000000000000000000000000000011;
	
	//x = 32'b10111111100100000000000000000000; //-1.125
	//y = 32'b01000000110000100000000000000000; //6.0625
	//r = 11000000110110100100000000000000 = -6.8203125
end
endmodule